`ifndef APB_MASTER_PKG_SV
`define APB_MASTER_PKG_SV

    `include "APB_master_seq_item.sv"
    `include "APB_master_sequences.sv"
    `include "APB_master_driver.sv"
    `include "APB_master_monitor.sv"
    `include "APB_master_sequencer.sv"
    `include "APB_master_agent.sv"

`endif // APB_MASTER_PKG_SV