package APB_env_pkg;

    import  uvm_pkg::*;
    import shared_pkg::*;

    `include "APB_config.sv"
    `include "APB_master_pkg.sv"
    `include "APB_slave_pkg.sv"
    `include "APB_coverage_collector.sv"
    `include "APB_scoreboard.sv"
    `include "APB_env.sv"

endpackage : APB_env_pkg