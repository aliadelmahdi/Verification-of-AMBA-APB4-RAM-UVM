
package APB_test_pkg;

    import  uvm_pkg::*;
    import  shared_pkg::*;
    import  APB_env_pkg::*;
    
    `include "APB_test_base.sv"

endpackage : APB_test_pkg