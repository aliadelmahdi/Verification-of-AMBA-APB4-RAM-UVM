`ifndef APB_MASTER_SEQUENCES_SV
`define APB_MASTER_SEQUENCES_SV

    `include "APB_master_reset_sequence.sv"
    `include "APB_master_main_sequence.sv"

`endif // APB_MASTER_SEQUENCES_SV
