`ifndef APB_SLAVE_SEQUENCES_SV
`define APB_SLAVE_SEQUENCES_SV

    `include "APB_slave_main_sequence.sv"

`endif // APB_SLAVE_SEQUENCES_SV